2
95 96 92 88 93 r 19 24 33 41 h 15 B 22 H 34 T
100 100 100 100 100 r 32 27 31 39 44 40 h 20 B 32 H 27 H
96 97 95 92 95 r 30 21 18 h 13 B 25 T
0 0 0 0 0 r h 37 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
4
